//--------------------------------------------------------------------------------
// File         : displaying.v
// Dependencies : 
// Description  : Demonstration of System Taks used for Displaying
//--------------------------------------------------------------------------------

module displaying();

  // $display is used to display data once, it and adds a newline character
  
  // $write is used to display data once, it doesnot add newline character
  
  // $strobe displays simulation data once at the end of current simulation time
  
  // $monitor displays data whenever it changes
  // $monitoroff can be used to disable monitoring for fast simulation
  // $monitoron can be used to enable monitoring

endmodule